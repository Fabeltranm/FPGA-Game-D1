module microfono
(
	input     Enable,
	input    [31:0]  data,
	output     Clk,
	output     ws,
	output     Dataout,
	output     Done,

);

endmodule
