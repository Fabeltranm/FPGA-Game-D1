﻿module	divisorFrec
(
	input           clkIn,
	output          clkOut
);
 endmodule
