module Ultrasonido	(

				output [0:7]	d,
				output 		trigg,
				output 		DONE,
				input 		ENABLE,
				input 		ECHO,
				input		clk

			 );


endmodule
