module touchScreen (input )