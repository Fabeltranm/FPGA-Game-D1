module Lectura	(

				output 		DONE,
				output	[7:0]	data,
				input		CLKOUT,
				input 		Rx

			 );


endmodule
