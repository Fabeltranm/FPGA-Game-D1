module contador		(
				
				output	[0:7] count,
				output	trigg,
				output	doneC
				input	ECHO,
				input	ENABLE
				
			);


endmodule
