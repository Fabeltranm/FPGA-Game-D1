module touchscreen #(
	parameter coordinate_x = 0,
	parameter coordinate_y = 0,
         
)(input init, input signal, input pulse, output coordinates);
