module Ultrasonido	(

				output Ren
				output R
				output Rm
				input f
				input Tro


			 );















endmodule
