module audio
(
	input             CLK,
	input      [15:0] D_IN,
	output            BCLK,
	output            LRCLK,
	output            DONE,
	output     	  D_OUT,

);
endmodule
