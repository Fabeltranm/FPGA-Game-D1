module	ultrasound
(
	input           clk,
	input           enable,
	input		echo,
	output   [7:0]  d,
	output		done,
	output          trigg
);
