module Touch	(

				output 		SDA,
				input 		SCL

			 );


endmodule
