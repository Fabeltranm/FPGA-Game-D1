module LVDS(CLK, Image, DataEnable, Channel0, Channel1, Channel2)
	( 
	input CLK,
	input Image,
	input DataEnable,
	output CLK,	
	output Channel0,
	output Channel1,
	output Channel2,
	);
	end
endmodule
