module microfono
(
	input     Enable,
	input    [31:0]  data,
	output     Clk,
	output     ws,
	output     Dataout,
	output     Done,
	parameter   count  = 0,

);

endmodule
