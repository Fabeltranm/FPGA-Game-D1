module microfono
(
	input     ws,
	output    [7:0]  Adress,
	input     Clk1,
	input     Reset,
	output     Done,
	output    [17:0]  Dataout
	input     data,
	input     select,
	output     Clk2,	

);

endmodule
