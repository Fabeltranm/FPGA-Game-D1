module Ultrasonido	(

				output [0:8]	d,
				output 		trigg,
				output 		DONE,
				input 		ENABLE,
				input 		ECHO,
				input		clk

			 );


endmodule
