﻿module	generadorPulsos
(
	input           clk,
	input		ECHO,
	input		enableP
	output          trigg,
	output		doneP,
	output	[7:0]	count
);
 endmodule
