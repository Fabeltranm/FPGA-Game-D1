module Touch	(

	output 		data,
	output		DONE,
	input		clk,
	input 		Rx
);


endmodule
