module	ultrasound
(
	input           clk,
	input           init,
	input		echo,
	output   [7:0]  d,
	output		done,
	output          trigg
);
