﻿module	divisorFrec	(
				input           CLKIN,
				output          CLKOUT
			);
endmodule
