module LVDS
	( 
	input CLK,
	input R,
	input G,
	input B,
	input DataEnable,
	output Channel 0,
	output Channel 1,
	output Channel 2,
	output CLK,
	);
endmodule
