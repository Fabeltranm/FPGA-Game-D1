module contador		(
				
				output	[7:0] count,
				output	trigg,
				output	calculate,
				input	ECHO,
				input	ENABLE,
				input	CLKOUT
				
			);


endmodule
