module Touch	(

	output 		data,
	output		DONE,
	output		clk,
	input 		Rx
);


endmodule
