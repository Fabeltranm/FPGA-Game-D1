module contador		(
				
				output	[7:0] count,
				output	trigg,
				output	doneC,
				input	ECHO,
				input	ENABLE,
				input	CLKOUT
				
			);


endmodule
