module microfono
(
	input     bclk,
	output    [7:0]  Adress,
	input     sdmode,
	input     Reset,
	input     [14:0]  Datain,
	input     select,
	output    done,	

);

endmodule
