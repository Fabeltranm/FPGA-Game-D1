module	multiplo	(
				input   [7:0]   count,
				input		calculate,
				output		DONE,
				output	[7:0]	d
			);
endmodule
