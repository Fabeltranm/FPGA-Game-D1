module Ultrasonido	(

				output Ren,
				output [0:8] R,
				output Rm,
				output i,
				input f,
				input Tro


			 );



endmodule
