module	divisorfrec	(
				input           clk,
				output          CLKOUT
			);
endmodule
