module proyecto
	( 
	input [15:0] dataIN,
	input EN,
	input reset,
	input CLK
	input MISO,
	input RW,
	input [15:0] addres,
	output [15:0] dataOUT,
	output DONE,
	output MOSI,
	output CS,
	);






endmodule
