module proyecto
	( 
	input [15:0] dataIN,
	input EN,
	input reset,
	input CLK
	input DATA0,
	input RW,
	input [7:0] addres,
	output [15:0] dataOUT,
	output DONE,
	output CMD,
	output DATA3,
	);






endmodule
