﻿module	generadorPulsos
(
	input		ECHO,
	output          trigg
);
 endmodule
