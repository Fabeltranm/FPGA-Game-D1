module LVDS
	( 
	input CLK,
	input Image,
	input DataEnable,
	output Channel 0,
	output Channel 1,
	output Channel 2,
	);
endmodule
