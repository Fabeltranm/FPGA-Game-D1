module Touch	(

				output 		SDA1,
				input		SDA2,
				input 		SCL

			 );


endmodule
