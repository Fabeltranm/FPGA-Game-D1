﻿module	divisor
(
	input           count,
	input		enable
	output		done,
	output	[7:0]	d
);